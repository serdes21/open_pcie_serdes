************************************************************************
* auCdl Netlist:
* 
* Library Name:  SerDes_16G_NRZ
* Top Cell Name: Half_rate_NRZ_16G
* View Name:     schematic
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    C2MOS_Latch
* View Name:    schematic
************************************************************************

.SUBCKT C2MOS_Latch AVDD AVSS CLK DO DO_B VO VO_B
*.PININFO CLK:I DO:I DO_B:I VO:O VO_B:O AVDD:B AVSS:B
MNM6 VO net079 AVSS AVSS N_1P05_HLPELVT W=400n L=30n M=3
MNM9 VO_B net078 AVSS AVSS N_1P05_HLPELVT W=400n L=30n M=3
MNM7 net079 net073 AVSS AVSS N_1P05_HLPELVT W=400n L=30n M=1
MNM8 net078 net072 AVSS AVSS N_1P05_HLPELVT W=400n L=30n M=1
MNM2 net073 DO_B net049 AVSS N_1P05_HLPELVT W=1.5u L=30n M=1
MNM10 net072 net073 AVSS AVSS N_1P05_HLPELVT W=500n L=30n M=1
MNM1 net049 CLKI AVSS AVSS N_1P05_HLPELVT W=1.5u L=30n M=1
MNM5 net073 net072 AVSS AVSS N_1P05_HLPELVT W=500n L=30n M=1
MNM0 net072 DO net049 AVSS N_1P05_HLPELVT W=1.5u L=30n M=1
MNM4 CLKI CLK AVSS AVSS N_1P05_HLPELVT W=100n L=30n M=1
MNM3 CLK AVDD CLKT AVSS N_1P05_HLPELVT W=100n L=30n M=1
MPM6 VO net079 AVDD AVDD P_1P05_HLPELVT W=600n L=30n M=3
MPM9 VO_B net078 AVDD AVDD P_1P05_HLPELVT W=600n L=30n M=3
MPM7 net079 net073 AVDD AVDD P_1P05_HLPELVT W=600n L=30n M=1
MPM8 net078 net072 AVDD AVDD P_1P05_HLPELVT W=600n L=30n M=1
MPM0 net073 DO_B net050 AVDD P_1P05_HLPELVT W=2.4u L=30n M=1
MPM10 net072 net073 AVDD AVDD P_1P05_HLPELVT W=900n L=30n M=1
MPM1 net050 CLKT AVDD AVDD P_1P05_HLPELVT W=4.8u L=30n M=1
MPM5 net073 net072 AVDD AVDD P_1P05_HLPELVT W=900n L=30n M=1
MPM3 net072 DO net050 AVDD P_1P05_HLPELVT W=2.4u L=30n M=1
MPM4 CLKI CLK AVDD AVDD P_1P05_HLPELVT W=230n L=30n M=1
MPM2 CLK AVSS CLKT AVDD P_1P05_HLPELVT W=230n L=30n M=1
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    INV_2
* View Name:    schematic
************************************************************************

.SUBCKT INV_2 AVDD AVSS CK CKB CLK
*.PININFO CLK:I CK:O CKB:O AVDD:B AVSS:B
MPM0 CK CKB AVDD AVDD P_1P05_HLPELVT W=900n L=30n M=8
MPM8 CKB CLK AVDD AVDD P_1P05_HLPELVT W=900n L=30n M=4
MNM0 CK CKB AVSS AVSS N_1P05_HLPELVT W=500n L=30n M=8
MNM8 CKB CLK AVSS AVSS N_1P05_HLPELVT W=500n L=30n M=4
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    High_speed_pre_driver
* View Name:    schematic
************************************************************************

.SUBCKT High_speed_pre_driver AVDD AVSS VIN VOUT
*.PININFO VIN:I VOUT:O AVDD:B AVSS:B
MPM15 VOUT net58 AVDD AVDD P_1P05_HLPELVT W=128u L=30n M=1
MPM1 net58 net57 AVDD AVDD P_1P05_HLPELVT W=64u L=30n M=1
MPM10 net57 net56 AVDD AVDD P_1P05_HLPELVT W=32u L=30n M=1
MPM8 net56 net55 AVDD AVDD P_1P05_HLPELVT W=16u L=30n M=1
MPM0 net55 VIN AVDD AVDD P_1P05_HLPELVT W=8u L=30n M=1
MNM16 VOUT net58 AVSS AVSS N_1P05_HLPELVT W=64u L=30n M=1
MNM1 net58 net57 AVSS AVSS N_1P05_HLPELVT W=32u L=30n M=1
MNM11 net57 net56 AVSS AVSS N_1P05_HLPELVT W=16u L=30n M=1
MNM10 net56 net55 AVSS AVSS N_1P05_HLPELVT W=8u L=30n M=1
MNM0 net55 VIN AVSS AVSS N_1P05_HLPELVT W=4u L=30n M=1
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    High_Speed_MUX_2_1
* View Name:    schematic
************************************************************************

.SUBCKT High_Speed_MUX_2_1 AVDD AVSS CLK D0 D1 VOUT
*.PININFO CLK:I D0:I D1:I VOUT:O AVDD:B AVSS:B
MNM17 VOUT net107 AVSS AVSS N_1P05_HLPELVT W=300n L=30n M=8
MNM16 net107 net106 AVSS AVSS N_1P05_HLPELVT W=300n L=30n M=4
MNM15 net106 OUT AVSS AVSS N_1P05_HLPELVT W=300n L=30n M=2
MNM14 OUT CLKT net109 AVSS N_1P05_HLPELVT W=300n L=30n M=1
MNM13 net109 D1 AVSS AVSS N_1P05_HLPELVT W=1u L=30n M=2
MNM12 OUT CLKI net111 AVSS N_1P05_HLPELVT W=300n L=30n M=1
MNM11 net111 D0 AVSS AVSS N_1P05_HLPELVT W=1u L=30n M=2
MNM10 CLKI CLK AVSS AVSS N_1P05_HLPELVT W=100n L=30n M=1
MNM9 CLK AVDD CLKT AVSS N_1P05_HLPELVT W=100n L=30n M=1
MPM17 VOUT net107 AVDD AVDD P_1P05_HLPELVT W=500n L=30n M=8
MPM16 net107 net106 AVDD AVDD P_1P05_HLPELVT W=500n L=30n M=4
MPM15 net106 OUT AVDD AVDD P_1P05_HLPELVT W=500n L=30n M=2
MPM14 net108 D1 AVDD AVDD P_1P05_HLPELVT W=1.2u L=30n M=2
MPM13 OUT CLKI net108 AVDD P_1P05_HLPELVT W=400n L=30n M=1
MPM12 net110 D0 AVDD AVDD P_1P05_HLPELVT W=1.2u L=30n M=2
MPM11 OUT CLKT net110 AVDD P_1P05_HLPELVT W=400n L=30n M=1
MPM10 CLKI CLK AVDD AVDD P_1P05_HLPELVT W=230n L=30n M=1
MPM8 CLK AVSS CLKT AVDD P_1P05_HLPELVT W=230n L=30n M=1
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    CML_pmos
* View Name:    schematic
************************************************************************

.SUBCKT CML_pmos AVDD AVSS MN<0> MN<1> MN<2> MP<0> MP<1> MP<2> VREF on op
*.PININFO MN<0>:I MN<1>:I MN<2>:I MP<0>:I MP<1>:I MP<2>:I VREF:I on:O op:O 
*.PININFO AVDD:B AVSS:B
MPM7 on MN<2> net8 AVDD P_1P05_HLPELVT W=15u L=30n M=1
MPM6 net8 AVDD AVDD AVDD P_1P05_HLPELVT W=37.5u L=30n M=1
MPM8 op MP<2> net8 AVDD P_1P05_HLPELVT W=15u L=30n M=1
MPM2 op MN<1> net6 AVDD P_1P05_HLPELVT W=60.2u L=30n M=1
MPM0 net6 VREF AVDD AVDD P_1P05_HLPELVT W=150.8u L=30n M=1
MPM1 on MP<1> net6 AVDD P_1P05_HLPELVT W=60.2u L=30n M=1
MPM4 on MN<0> net3 AVDD P_1P05_HLPELVT W=6.7u L=30n M=1
MPM3 op MP<0> net3 AVDD P_1P05_HLPELVT W=6.7u L=30n M=1
MPM5 net3 AVDD AVDD AVDD P_1P05_HLPELVT W=16.8u L=30n M=1
RR24 AVSS op 49.8601 $SUB=AVSS $[RNNPO_HLP] $W=4.8u $L=900n M=1
RR25 AVSS on 49.8601 $SUB=AVSS $[RNNPO_HLP] $W=4.8u $L=900n M=1
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    PLatch_TG
* View Name:    schematic
************************************************************************

.SUBCKT PLatch_TG AVDD AVSS CLK D Q
*.PININFO CLK:I D:I Q:O AVDD:B AVSS:B
MNM5 CLKI CLK AVSS AVSS N_1P05_HLPELVT W=100n L=30n M=1
MNM4 Q DIT AVSS AVSS N_1P05_HLPELVT W=100n L=30n M=2
MNM3 DI CLKT DIT AVSS N_1P05_HLPELVT W=100n L=30n M=2
MNM2 QI CLKI DIT AVSS N_1P05_HLPELVT W=100n L=30n M=2
MNM1 QI Q AVSS AVSS N_1P05_HLPELVT W=100n L=30n M=2
MNM0 DI D AVSS AVSS N_1P05_HLPELVT W=100n L=30n M=2
MNM6 CLK AVDD CLKT AVSS N_1P05_HLPELVT W=100n L=30n M=1
MPM5 CLKI CLK AVDD AVDD P_1P05_HLPELVT W=230n L=30n M=1
MPM4 Q DIT AVDD AVDD P_1P05_HLPELVT W=230n L=30n M=2
MPM3 DI CLKI DIT AVDD P_1P05_HLPELVT W=230n L=30n M=2
MPM2 QI CLKT DIT AVDD P_1P05_HLPELVT W=230n L=30n M=2
MPM1 QI Q AVDD AVDD P_1P05_HLPELVT W=230n L=30n M=2
MPM0 DI D AVDD AVDD P_1P05_HLPELVT W=230n L=30n M=2
MPM6 CLK AVSS CLKT AVDD P_1P05_HLPELVT W=230n L=30n M=1
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    DFF_C2mos_td
* View Name:    schematic
************************************************************************

.SUBCKT DFF_C2mos_td AVDD AVSS CLK D Q
*.PININFO CLK:I D:I Q:O AVDD:B AVSS:B
MPM6 CLK AVSS CLKT AVDD P_1P05_HLPELVT W=230n L=30n M=1
MPM4 Q net43 AVDD AVDD P_1P05_HLPELVT W=500n L=30n M=4
MPM8 net43 Qt AVDD AVDD P_1P05_HLPELVT W=500n L=30n M=1
MPM3 Qt CLKT net44 AVDD P_1P05_HLPELVT W=230n L=30n M=1
MPM2 net44 D1 AVDD AVDD P_1P05_HLPELVT W=400n L=30n M=1
MPM1 D1 CLKI net46 AVDD P_1P05_HLPELVT W=230n L=30n M=1
MPM5 CLKI CLK AVDD AVDD P_1P05_HLPELVT W=230n L=30n M=1
MPM0 net46 D AVDD AVDD P_1P05_HLPELVT W=400n L=30n M=1
MNM5 CLKI CLK AVSS AVSS N_1P05_HLPELVT W=100n L=30n M=1
MNM4 Q net43 AVSS AVSS N_1P05_HLPELVT W=300n L=30n M=4
MNM8 net43 Qt AVSS AVSS N_1P05_HLPELVT W=300n L=30n M=1
MNM2 Qt CLKI net45 AVSS N_1P05_HLPELVT W=200n L=30n M=1
MNM3 net45 D1 AVSS AVSS N_1P05_HLPELVT W=200n L=30n M=1
MNM6 CLK AVDD CLKT AVSS N_1P05_HLPELVT W=100n L=30n M=1
MNM0 D1 CLKT net47 AVSS N_1P05_HLPELVT W=200n L=30n M=1
MNM1 net47 D AVSS AVSS N_1P05_HLPELVT W=200n L=30n M=1
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    SEL2_1_TG
* View Name:    schematic
************************************************************************

.SUBCKT SEL2_1_TG AVDD AVSS CLK D1 D2 Q
*.PININFO CLK:I D1:I D2:I Q:O AVDD:B AVSS:B
MNM5 CLKI CLK AVSS AVSS N_1P05_HLPELVT W=100n L=30n M=1
MNM3 Q net64 AVSS AVSS N_1P05_HLPELVT W=300n L=30n M=4
MNM2 net64 DQ AVSS AVSS N_1P05_HLPELVT W=300n L=30n M=1
MNM1 D2 CLKT DQ AVSS N_1P05_HLPELVT W=200n L=30n M=1
MNM0 D1 CLKI DQ AVSS N_1P05_HLPELVT W=200n L=30n M=1
MNM6 CLK AVDD CLKT AVSS N_1P05_HLPELVT W=100n L=30n M=1
MPM5 CLKI CLK AVDD AVDD P_1P05_HLPELVT W=230n L=30n M=1
MPM3 Q net64 AVDD AVDD P_1P05_HLPELVT W=500n L=30n M=4
MPM2 net64 DQ AVDD AVDD P_1P05_HLPELVT W=500n L=30n M=1
MPM1 D2 CLKI DQ AVDD P_1P05_HLPELVT W=400n L=30n M=1
MPM0 D1 CLKT DQ AVDD P_1P05_HLPELVT W=400n L=30n M=1
MPM6 CLK AVSS CLKT AVDD P_1P05_HLPELVT W=230n L=30n M=1
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    5Latch_MUX2_1_TG
* View Name:    schematic
************************************************************************

.SUBCKT 5Latch_MUX2_1_TG AVDD AVSS CK_0 CK_90 D1 D2 Q
*.PININFO CK_0:I CK_90:I D1:I D2:I Q:O AVDD:B AVSS:B
Xi2 AVDD AVSS CK_0 net28 D2_d2 / PLatch_TG
Xi0 AVDD AVSS CK_0 D1 D1_d1 / DFF_C2mos_td
Xi1 AVDD AVSS CK_0 D2 net28 / DFF_C2mos_td
Xi3 AVDD AVSS CK_90 D1_d1 D2_d2 Q / SEL2_1_TG
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    Serial32_2__buffer
* View Name:    schematic
************************************************************************

.SUBCKT Serial32_2__buffer AVDD AVSS D DI DT
*.PININFO D:I DI:O DT:O AVDD:B AVSS:B
MNM2 DI net57 AVSS AVSS N_1P05_HLPELVT W=300n L=30n M=4
MNM0 DT net55 AVSS AVSS N_1P05_HLPELVT W=300n L=30n M=4
MNM8 net55 D AVSS AVSS N_1P05_HLPELVT W=300n L=30n M=1
MNM1 D AVDD net57 AVSS N_1P05_HLPELVT W=300n L=30n M=1
MPM2 DI net57 AVDD AVDD P_1P05_HLPELVT W=500n L=30n M=4
MPM0 DT net55 AVDD AVDD P_1P05_HLPELVT W=500n L=30n M=4
MPM8 net55 D AVDD AVDD P_1P05_HLPELVT W=500n L=30n M=1
MPM1 D AVSS net57 AVDD P_1P05_HLPELVT W=500n L=30n M=1
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    3Latch_MUX2_1_TG
* View Name:    schematic
************************************************************************

.SUBCKT 3Latch_MUX2_1_TG AVDD AVSS CK_0 CK_90 D1 D2 Q
*.PININFO CK_0:I CK_90:I D1:I D2:I Q:O AVDD:B AVSS:B
Xi1 AVDD AVSS CK_0 D1 D1_d1 / DFF_C2mos_td
Xi2 AVDD AVSS CK_90 D1_d1 D2_d2 Q / SEL2_1_TG
Xi0 AVDD AVSS CK_0 D2 D2_d2 / PLatch_TG
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    Serial32_2__Tree_MUX2_1_TG
* View Name:    schematic
************************************************************************

.SUBCKT Serial32_2__Tree_MUX2_1_TG AVDD AVSS CK16_0 CK16_90 CK32_0 CK32_90 
+ CK4_0 CK4_90 CK8_0 CK8_90 D2I<0> D2I<1> D2T<0> D2T<1> D32<0> D32<10> D32<11> 
+ D32<12> D32<13> D32<14> D32<15> D32<16> D32<17> D32<18> D32<19> D32<1> 
+ D32<20> D32<21> D32<22> D32<23> D32<24> D32<25> D32<26> D32<27> D32<28> 
+ D32<29> D32<2> D32<30> D32<31> D32<3> D32<4> D32<5> D32<6> D32<7> D32<8> 
+ D32<9>
*.PININFO CK4_0:I CK4_90:I CK8_0:I CK8_90:I CK16_0:I CK16_90:I CK32_0:I 
*.PININFO CK32_90:I D32<0>:I D32<1>:I D32<2>:I D32<3>:I D32<4>:I D32<5>:I 
*.PININFO D32<6>:I D32<7>:I D32<8>:I D32<9>:I D32<10>:I D32<11>:I D32<12>:I 
*.PININFO D32<13>:I D32<14>:I D32<15>:I D32<16>:I D32<17>:I D32<18>:I 
*.PININFO D32<19>:I D32<20>:I D32<21>:I D32<22>:I D32<23>:I D32<24>:I 
*.PININFO D32<25>:I D32<26>:I D32<27>:I D32<28>:I D32<29>:I D32<30>:I 
*.PININFO D32<31>:I D2I<0>:O D2I<1>:O D2T<0>:O D2T<1>:O AVDD:B AVSS:B
Xi0 AVDD AVSS CK32_0 CK32_90 D32<0> D32<16> D16<0> / 5Latch_MUX2_1_TG
Xi15 AVDD AVSS CK32_0 CK32_90 D32<8> D32<24> D16<8> / 5Latch_MUX2_1_TG
Xi14 AVDD AVSS CK32_0 CK32_90 D32<9> D32<25> D16<9> / 5Latch_MUX2_1_TG
Xi1 AVDD AVSS CK32_0 CK32_90 D32<1> D32<17> D16<1> / 5Latch_MUX2_1_TG
Xi13 AVDD AVSS CK32_0 CK32_90 D32<10> D32<26> D16<10> / 5Latch_MUX2_1_TG
Xi2 AVDD AVSS CK32_0 CK32_90 D32<2> D32<18> D16<2> / 5Latch_MUX2_1_TG
Xi7 AVDD AVSS CK32_0 CK32_90 D32<7> D32<23> D16<7> / 5Latch_MUX2_1_TG
Xi3 AVDD AVSS CK32_0 CK32_90 D32<3> D32<19> D16<3> / 5Latch_MUX2_1_TG
Xi12 AVDD AVSS CK32_0 CK32_90 D32<11> D32<27> D16<11> / 5Latch_MUX2_1_TG
Xi11 AVDD AVSS CK32_0 CK32_90 D32<12> D32<28> D16<12> / 5Latch_MUX2_1_TG
Xi10 AVDD AVSS CK32_0 CK32_90 D32<13> D32<29> D16<13> / 5Latch_MUX2_1_TG
Xi5 AVDD AVSS CK32_0 CK32_90 D32<5> D32<21> D16<5> / 5Latch_MUX2_1_TG
Xi9 AVDD AVSS CK32_0 CK32_90 D32<14> D32<30> D16<14> / 5Latch_MUX2_1_TG
Xi6 AVDD AVSS CK32_0 CK32_90 D32<6> D32<22> D16<6> / 5Latch_MUX2_1_TG
Xi8 AVDD AVSS CK32_0 CK32_90 D32<15> D32<31> D16<15> / 5Latch_MUX2_1_TG
Xi4 AVDD AVSS CK32_0 CK32_90 D32<4> D32<20> D16<4> / 5Latch_MUX2_1_TG
Xi28 AVDD AVSS D2<0> D2I<0> D2T<0> / Serial32_2__buffer
Xi29 AVDD AVSS D2<1> D2I<1> D2T<1> / Serial32_2__buffer
Xi33 AVDD AVSS CK4_0 CK4_90 D4<0> D4<2> D2<0> / 3Latch_MUX2_1_TG
Xi32 AVDD AVSS CK4_0 CK4_90 D4<1> D4<3> D2<1> / 3Latch_MUX2_1_TG
Xi24 AVDD AVSS CK8_0 CK8_90 D8<0> D8<4> D4<0> / 3Latch_MUX2_1_TG
Xi16 AVDD AVSS CK16_0 CK16_90 D16<0> D16<8> D8<0> / 3Latch_MUX2_1_TG
Xi25 AVDD AVSS CK8_0 CK8_90 D8<1> D8<5> D4<1> / 3Latch_MUX2_1_TG
Xi17 AVDD AVSS CK16_0 CK16_90 D16<1> D16<9> D8<1> / 3Latch_MUX2_1_TG
Xi26 AVDD AVSS CK8_0 CK8_90 D8<2> D8<6> D4<2> / 3Latch_MUX2_1_TG
Xi18 AVDD AVSS CK16_0 CK16_90 D16<2> D16<10> D8<2> / 3Latch_MUX2_1_TG
Xi23 AVDD AVSS CK16_0 CK16_90 D16<7> D16<15> D8<7> / 3Latch_MUX2_1_TG
Xi27 AVDD AVSS CK8_0 CK8_90 D8<3> D8<7> D4<3> / 3Latch_MUX2_1_TG
Xi19 AVDD AVSS CK16_0 CK16_90 D16<3> D16<11> D8<3> / 3Latch_MUX2_1_TG
Xi21 AVDD AVSS CK16_0 CK16_90 D16<5> D16<13> D8<5> / 3Latch_MUX2_1_TG
Xi22 AVDD AVSS CK16_0 CK16_90 D16<6> D16<14> D8<6> / 3Latch_MUX2_1_TG
Xi20 AVDD AVSS CK16_0 CK16_90 D16<4> D16<12> D8<4> / 3Latch_MUX2_1_TG
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    div_2_4_8
* View Name:    schematic
************************************************************************

.SUBCKT div_2_4_8 AVDD AVSS CLK EN Q
*.PININFO CLK:I EN:I Q:O AVDD:B AVSS:B
MPM14 Q net97 AVDD AVDD P_1P05_HLPELVT W=600n L=30n M=1
MPM11 net97 EN AVDD AVDD P_1P05_HLPELVT W=500n L=200n M=1
MPM15 net97 net115 AVDD AVDD P_1P05_HLPELVT W=250n L=30n M=2
MPM16 net115 net112 AVDD AVDD P_1P05_HLPELVT W=250n L=30n M=1
MPM2 net118 net97 AVDD AVDD P_1P05_HLPELVT W=250n L=30n M=1
MPM1 net109 net112 net118 AVDD P_1P05_HLPELVT W=300n L=30n M=1
MPM8 net112 EN AVDD AVDD P_1P05_HLPELVT W=500n L=200n M=1
MPM10 net112 ENB CLK AVDD P_1P05_HLPELVT W=230n L=30n M=1
MPM3 ENB EN AVDD AVDD P_1P05_HLPELVT W=230n L=30n M=1
MNM19 Q net97 AVSS AVSS N_1P05_HLPELVT W=250n L=30n M=1
MNM16 net116 net115 AVSS AVSS N_1P05_HLPELVT W=120n L=30n M=1
MNM17 net97 net112 net116 AVSS N_1P05_HLPELVT W=150n L=30n M=1
MNM18 net115 net109 net117 AVSS N_1P05_HLPELVT W=200n L=30n M=1
MNM15 net117 net112 AVSS AVSS N_1P05_HLPELVT W=180n L=30n M=1
MNM2 net109 net97 AVSS AVSS N_1P05_HLPELVT W=150n L=30n M=1
MNM1 net112 EN CLK AVSS N_1P05_HLPELVT W=100n L=30n M=1
MNM0 ENB EN AVSS AVSS N_1P05_HLPELVT W=100n L=30n M=1
.ENDS

************************************************************************
* Library Name: SerDes_16G_NRZ
* Cell Name:    Half_rate_NRZ_16G
* View Name:    schematic
************************************************************************

.SUBCKT Half_rate_NRZ_16G AVDD AVDD_1P2 AVSS CK_8G CK_B_8G D32<0> D32<10> 
+ D32<11> D32<12> D32<13> D32<14> D32<15> D32<16> D32<17> D32<18> D32<19> 
+ D32<1> D32<20> D32<21> D32<22> D32<23> D32<24> D32<25> D32<26> D32<27> 
+ D32<28> D32<29> D32<2> D32<30> D32<31> D32<3> D32<4> D32<5> D32<6> D32<7> 
+ D32<8> D32<9> EN ON OP VREF
*.PININFO CK_8G:I CK_B_8G:I D32<0>:I D32<1>:I D32<2>:I D32<3>:I D32<4>:I 
*.PININFO D32<5>:I D32<6>:I D32<7>:I D32<8>:I D32<9>:I D32<10>:I D32<11>:I 
*.PININFO D32<12>:I D32<13>:I D32<14>:I D32<15>:I D32<16>:I D32<17>:I 
*.PININFO D32<18>:I D32<19>:I D32<20>:I D32<21>:I D32<22>:I D32<23>:I 
*.PININFO D32<24>:I D32<25>:I D32<26>:I D32<27>:I D32<28>:I D32<29>:I 
*.PININFO D32<30>:I D32<31>:I EN:I VREF:I ON:O OP:O AVDD:B AVDD_1P2:B AVSS:B
Xi21 AVDD AVSS CK_8G D2T<0> D2I<0> net0111 net0112 / C2MOS_Latch
Xi39 AVDD AVSS CK_B_8G BN<1> BP<1> BN<2> BP<2> / C2MOS_Latch
Xi40 AVDD AVSS CK_8G BN<0> BP<0> BN<1> BP<1> / C2MOS_Latch
Xi41 AVDD AVSS CK_B_8G net0108 net0107 BN<0> BP<0> / C2MOS_Latch
Xi42 AVDD AVSS CK_8G D2T<1> D2I<1> net0108 net0107 / C2MOS_Latch
Xi26 AVDD AVSS CK_8G net0110 net0109 AN<0> AP<0> / C2MOS_Latch
Xi36 AVDD AVSS CK_B_8G AN<0> AP<0> AN<1> AP<1> / C2MOS_Latch
Xi38 AVDD AVSS CK_8G AN<1> AP<1> AN<2> AP<2> / C2MOS_Latch
Xi24 AVDD AVSS CK_B_8G net0111 net0112 net0110 net0109 / C2MOS_Latch
Xi22 AVDD AVSS CK_2G CK_B_2G CK1_2G / INV_2
Xi23 AVDD AVSS CK_1G CK_B_1G CK1_1G / INV_2
Xi16 AVDD AVSS CK_4G CK_B_4G CK1_4G / INV_2
Xi14 AVDD AVSS CK_0P5G CK_B_0P5G CK1_0P5G / INV_2
Xi5 AVDD AVSS MN<0> MMN<0> / High_speed_pre_driver
Xi4 AVDD AVSS MP<0> MMP<0> / High_speed_pre_driver
Xi8 AVDD AVSS MP<1> MMP<1> / High_speed_pre_driver
Xi6 AVDD AVSS MN<1> MMN<1> / High_speed_pre_driver
Xi10 AVDD AVSS MN<2> MMN<2> / High_speed_pre_driver
Xi12 AVDD AVSS MP<2> MMP<2> / High_speed_pre_driver
Xi17 AVDD AVSS CK_8G AN<0> BN<0> MN<0> / High_Speed_MUX_2_1
Xi27 AVDD AVSS CK_8G AN<2> BN<2> MN<2> / High_Speed_MUX_2_1
Xi28 AVDD AVSS CK_B_8G AN<1> BN<1> MN<1> / High_Speed_MUX_2_1
Xi18 AVDD AVSS CK_8G AP<0> BP<0> MP<0> / High_Speed_MUX_2_1
Xi19 AVDD AVSS CK_B_8G AP<1> BP<1> MP<1> / High_Speed_MUX_2_1
Xi20 AVDD AVSS CK_8G AP<2> BP<2> MP<2> / High_Speed_MUX_2_1
Xi0 AVDD_1P2 AVSS MMN<0> MMN<1> MMN<2> MMP<0> MMP<1> MMP<2> VREF ON OP / 
+ CML_pmos
XI1 AVDD AVSS CK_1G CK_B_1G CK_0P5G CK_B_0P5G CK_4G CK_B_4G CK_2G CK_B_2G 
+ D2I<0> D2I<1> D2T<0> D2T<1> D32<0> D32<10> D32<11> D32<12> D32<13> D32<14> 
+ D32<15> D32<16> D32<17> D32<18> D32<19> D32<1> D32<20> D32<21> D32<22> 
+ D32<23> D32<24> D32<25> D32<26> D32<27> D32<28> D32<29> D32<2> D32<30> 
+ D32<31> D32<3> D32<4> D32<5> D32<6> D32<7> D32<8> D32<9> / 
+ Serial32_2__Tree_MUX2_1_TG
Xi3 AVDD AVSS CK_8G EN CK1_4G / div_2_4_8
Xi1 AVDD AVSS CK_2G EN CK1_1G / div_2_4_8
Xi2 AVDD AVSS CK_4G EN CK1_2G / div_2_4_8
Xi15 AVDD AVSS CK_1G EN CK1_0P5G / div_2_4_8
.ENDS

